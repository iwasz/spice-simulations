*******************************************************************
* Model name       : 1N5817
* Description      : Low Drop Power Schottky Diode
* Package type     : DO-41
*******************************************************************
.MODEL 1N5817 D IS=698.22E-9 N=1.0015 RS=35.457E-3 IKF=6.0924 CJO=345.48E-12
+ M=.45399 VJ=.3905 ISR=2.0219E-6 NR=4.9950 EG=.69 XTI=2 TT=0 FC=0.5
*$

